module main;

    initial begin
        $display("Icarus Verilog is working!");
        $finish;
    end

endmodule

